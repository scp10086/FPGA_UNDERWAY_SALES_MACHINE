----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 2019/09/05 15:55:52
-- Design Name: 
-- Module Name: choose_price - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.All;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity choose_price is
  Port (clk,switch4,switch5,switch6,switch7,confirm:in std_logic; --���ĸ����طֱ��Ӧ�ſ���ѡƱ�ۣ�2Ԫ��3Ԫ��5Ԫ��7Ԫ
        --led4,led5,led6,led7:out std_logic;
        dispdata :out std_logic_vector(31 downto 0);
        get_present_state:in std_logic_vector(3 downto 0);
        ticket_price:out std_logic_vector(3 downto 0);
        flag0:out std_logic);
end choose_price;

architecture Behavioral of choose_price is


signal confirm0,switch40,switch50,switch60,switch70:std_logic;
begin

process(clk)
begin
if (clk'event and clk='1') then
    confirm0<=confirm;
    switch40<=switch4;
    switch50<=switch5;
    switch60<=switch6;
    switch70<=switch7;
end if;
end process;

process(clk,confirm,switch4,switch5,switch6,switch7,get_present_state)
begin
  if (clk'event and clk='1') then
  
  if(get_present_state="0011") then
  flag0<='1'; --���������ѡƱ��������� ��ô���־λΪ1
  
    if (switch4='1'and switch40='0') then 
       if(confirm='1'and confirm0='0') then ticket_price<="0010";dispdata<=x"00000002";end if;
    end if;
    
    if (switch5='1'and switch50='0') then 
       if(confirm='1'and confirm0='0') then ticket_price<="0011";dispdata<=x"00000003";end if;
    end if;

    if (switch6='1'and switch60='0') then 
       if(confirm='1'and confirm0='0') then ticket_price<="0101";dispdata<=x"00000005";end if;
    end if;
    
    if (switch7='1'and switch70='0') then 
           if(confirm='1'and confirm0='0') then ticket_price<="0111";dispdata<=x"00000007";end if;
        end if;

  end if;
  else flag0<='0';
end if;
end process;

end Behavioral;
